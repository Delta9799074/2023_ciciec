/*
Copyright (c) 2019 Alibaba Group Holding Limited

Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software is furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

*/
module retu_top(
  hmain0_ismc_s0_haddr,
  hmain0_ismc_s0_hprot,
  hmain0_ismc_s0_hsel,
  hmain0_ismc_s0_hsize,
  hmain0_ismc_s0_htrans,
  hmain0_ismc_s0_hwdata,
  hmain0_ismc_s0_hwrite,
  hmain0_smc_s2_haddr,
  hmain0_smc_s2_hprot,
  hmain0_smc_s2_hsel,
  hmain0_smc_s2_hsize,
  hmain0_smc_s2_htrans,
  hmain0_smc_s2_hwdata,
  hmain0_smc_s2_hwrite,
  hmain0_smc_s3_haddr,
  hmain0_smc_s3_hprot,
  hmain0_smc_s3_hsel,
  hmain0_smc_s3_hsize,
  hmain0_smc_s3_htrans,
  hmain0_smc_s3_hwdata,
  hmain0_smc_s3_hwrite,
  hmain0_smc_s4_haddr,
  hmain0_smc_s4_hprot,
  hmain0_smc_s4_hsel,
  hmain0_smc_s4_hsize,
  hmain0_smc_s4_htrans,
  hmain0_smc_s4_hwdata,
  hmain0_smc_s4_hwrite,
  ismc_hmain0_s0_hrdata,
  ismc_hmain0_s0_hready,
  ismc_hmain0_s0_hresp,
  pmu_smc_hclk,
  pmu_smc_hrst_b,
  smc_hmain0_s2_hrdata,
  smc_hmain0_s2_hready,
  smc_hmain0_s2_hresp,
  smc_hmain0_s3_hrdata,
  smc_hmain0_s3_hready,
  smc_hmain0_s3_hresp,
  smc_hmain0_s4_hrdata,
  smc_hmain0_s4_hready,
  smc_hmain0_s4_hresp,

  //40个信号
hmain0_dummy3_s11_haddr,     
hmain0_dummy3_s11_hprot,    
hmain0_dummy3_s11_hsel,     
hmain0_dummy3_s11_hsize,    
hmain0_dummy3_s11_htrans,   
hmain0_dummy3_s11_hwdata,   
hmain0_dummy3_s11_hwrite, 
hmain0_dummy0_s7_haddr,     
hmain0_dummy0_s7_hprot,     
hmain0_dummy0_s7_hsel,      
hmain0_dummy0_s7_hsize,     
hmain0_dummy0_s7_htrans,    
hmain0_dummy0_s7_hwdata,    
hmain0_dummy0_s7_hwrite,    
hmain0_dummy1_s8_haddr,       
hmain0_dummy1_s8_hprot,     
hmain0_dummy1_s8_hsel,      
hmain0_dummy1_s8_hsize,     
hmain0_dummy1_s8_htrans,    
hmain0_dummy1_s8_hwdata,    
hmain0_dummy1_s8_hwrite,    
hmain0_dummy2_s9_haddr,       
hmain0_dummy2_s9_hprot,     
hmain0_dummy2_s9_hsel,      
hmain0_dummy2_s9_hsize,     
hmain0_dummy2_s9_htrans,    
hmain0_dummy2_s9_hwdata,    
hmain0_dummy2_s9_hwrite, 
dummy0_hmain0_s7_hrdata,    
dummy0_hmain0_s7_hready,    
dummy0_hmain0_s7_hresp,     
dummy1_hmain0_s8_hrdata,    
dummy1_hmain0_s8_hready,    
dummy1_hmain0_s8_hresp,     
dummy2_hmain0_s9_hrdata,    
dummy2_hmain0_s9_hready,    
dummy2_hmain0_s9_hresp,     
dummy3_hmain0_s11_hrdata,   
dummy3_hmain0_s11_hready,   
dummy3_hmain0_s11_hresp,

//1111
imemdummy0_hmain0_s1_hrdata, 
imemdummy0_hmain0_s1_hready, 
imemdummy0_hmain0_s1_hresp, 
hmain0_imemdummy0_s1_haddr, 
hmain0_imemdummy0_s1_hprot, 
hmain0_imemdummy0_s1_hsel,  
hmain0_imemdummy0_s1_hsize, 
hmain0_imemdummy0_s1_htrans, 
hmain0_imemdummy0_s1_hwdata, 
hmain0_imemdummy0_s1_hwrite

);
input   [31:0]  hmain0_ismc_s0_haddr; 
input   [3 :0]  hmain0_ismc_s0_hprot; 
input           hmain0_ismc_s0_hsel;  
input   [2 :0]  hmain0_ismc_s0_hsize; 
input   [1 :0]  hmain0_ismc_s0_htrans; 
input   [31:0]  hmain0_ismc_s0_hwdata; 
input           hmain0_ismc_s0_hwrite; 
input   [31:0]  hmain0_smc_s2_haddr;  
input   [3 :0]  hmain0_smc_s2_hprot;  
input           hmain0_smc_s2_hsel;   
input   [2 :0]  hmain0_smc_s2_hsize;  
input   [1 :0]  hmain0_smc_s2_htrans; 
input   [31:0]  hmain0_smc_s2_hwdata; 
input           hmain0_smc_s2_hwrite; 
input   [31:0]  hmain0_smc_s3_haddr;  
input   [3 :0]  hmain0_smc_s3_hprot;  
input           hmain0_smc_s3_hsel;   
input   [2 :0]  hmain0_smc_s3_hsize;  
input   [1 :0]  hmain0_smc_s3_htrans; 
input   [31:0]  hmain0_smc_s3_hwdata; 
input           hmain0_smc_s3_hwrite; 
input   [31:0]  hmain0_smc_s4_haddr;  
input   [3 :0]  hmain0_smc_s4_hprot;  
input           hmain0_smc_s4_hsel;   
input   [2 :0]  hmain0_smc_s4_hsize;  
input   [1 :0]  hmain0_smc_s4_htrans; 
input   [31:0]  hmain0_smc_s4_hwdata; 
input           hmain0_smc_s4_hwrite; 

input  [31:0]  hmain0_dummy3_s11_haddr;      
input  [3 :0]  hmain0_dummy3_s11_hprot;    
input          hmain0_dummy3_s11_hsel;     
input  [2 :0]  hmain0_dummy3_s11_hsize;    
input  [1 :0]  hmain0_dummy3_s11_htrans;   
input  [31:0]  hmain0_dummy3_s11_hwdata;   
input          hmain0_dummy3_s11_hwrite; 
input    [31:0]  hmain0_dummy0_s7_haddr;         
input    [3 :0]  hmain0_dummy0_s7_hprot;     
input            hmain0_dummy0_s7_hsel;      
input    [2 :0]  hmain0_dummy0_s7_hsize;     
input    [1 :0]  hmain0_dummy0_s7_htrans;    
input    [31:0]  hmain0_dummy0_s7_hwdata;    
input            hmain0_dummy0_s7_hwrite;    
input    [31:0]  hmain0_dummy1_s8_haddr;         
input    [3 :0]  hmain0_dummy1_s8_hprot;     
input            hmain0_dummy1_s8_hsel;      
input    [2 :0]  hmain0_dummy1_s8_hsize;     
input    [1 :0]  hmain0_dummy1_s8_htrans;    
input    [31:0]  hmain0_dummy1_s8_hwdata;    
input            hmain0_dummy1_s8_hwrite;    
input    [31:0]  hmain0_dummy2_s9_haddr;       
input    [3 :0]  hmain0_dummy2_s9_hprot;     
input            hmain0_dummy2_s9_hsel;      
input    [2 :0]  hmain0_dummy2_s9_hsize;     
input    [1 :0]  hmain0_dummy2_s9_htrans;    
input    [31:0]  hmain0_dummy2_s9_hwdata;    
input            hmain0_dummy2_s9_hwrite;

input    [31:0]  hmain0_imemdummy0_s1_haddr; 
input    [3 :0]  hmain0_imemdummy0_s1_hprot; 
input            hmain0_imemdummy0_s1_hsel;  
input    [2 :0]  hmain0_imemdummy0_s1_hsize; 
input    [1 :0]  hmain0_imemdummy0_s1_htrans; 
input    [31:0]  hmain0_imemdummy0_s1_hwdata; 
input            hmain0_imemdummy0_s1_hwrite;

input           pmu_smc_hclk;         
input           pmu_smc_hrst_b;     


output  [31:0]  ismc_hmain0_s0_hrdata; 
output          ismc_hmain0_s0_hready; 
output  [1 :0]  ismc_hmain0_s0_hresp; 
output  [31:0]  smc_hmain0_s2_hrdata; 
output          smc_hmain0_s2_hready; 
output  [1 :0]  smc_hmain0_s2_hresp;  
output  [31:0]  smc_hmain0_s3_hrdata; 
output          smc_hmain0_s3_hready; 
output  [1 :0]  smc_hmain0_s3_hresp;  
output  [31:0]  smc_hmain0_s4_hrdata; 
output          smc_hmain0_s4_hready; 
output  [1 :0]  smc_hmain0_s4_hresp;  

output    [31:0]  dummy3_hmain0_s11_hrdata;   
output            dummy3_hmain0_s11_hready;   
output    [1 :0]  dummy3_hmain0_s11_hresp; 
output    [31:0]  dummy0_hmain0_s7_hrdata;    
output            dummy0_hmain0_s7_hready;    
output    [1 :0]  dummy0_hmain0_s7_hresp;     
output    [31:0]  dummy1_hmain0_s8_hrdata;    
output            dummy1_hmain0_s8_hready;    
output    [1 :0]  dummy1_hmain0_s8_hresp;     
output    [31:0]  dummy2_hmain0_s9_hrdata;    
output            dummy2_hmain0_s9_hready;    
output    [1 :0]  dummy2_hmain0_s9_hresp;
//1111
output    [31:0]  imemdummy0_hmain0_s1_hrdata; 
output            imemdummy0_hmain0_s1_hready; 
output    [1 :0]  imemdummy0_hmain0_s1_hresp;

wire    [31:0]  hmain0_ismc_s0_haddr; 
wire    [3 :0]  hmain0_ismc_s0_hprot; 
wire            hmain0_ismc_s0_hsel;  
wire    [2 :0]  hmain0_ismc_s0_hsize; 
wire    [1 :0]  hmain0_ismc_s0_htrans; 
wire    [31:0]  hmain0_ismc_s0_hwdata; 
wire            hmain0_ismc_s0_hwrite; 
wire    [31:0]  hmain0_smc_s2_haddr;  
wire    [3 :0]  hmain0_smc_s2_hprot;  
wire            hmain0_smc_s2_hsel;   
wire    [2 :0]  hmain0_smc_s2_hsize;  
wire    [1 :0]  hmain0_smc_s2_htrans; 
wire    [31:0]  hmain0_smc_s2_hwdata; 
wire            hmain0_smc_s2_hwrite; 
wire    [31:0]  hmain0_smc_s3_haddr;  
wire    [3 :0]  hmain0_smc_s3_hprot;  
wire            hmain0_smc_s3_hsel;   
wire    [2 :0]  hmain0_smc_s3_hsize;  
wire    [1 :0]  hmain0_smc_s3_htrans; 
wire    [31:0]  hmain0_smc_s3_hwdata; 
wire            hmain0_smc_s3_hwrite; 
wire    [31:0]  hmain0_smc_s4_haddr;  
wire    [3 :0]  hmain0_smc_s4_hprot;  
wire            hmain0_smc_s4_hsel;   
wire    [2 :0]  hmain0_smc_s4_hsize;  
wire    [1 :0]  hmain0_smc_s4_htrans; 
wire    [31:0]  hmain0_smc_s4_hwdata; 
wire            hmain0_smc_s4_hwrite; 
wire    [31:0]  ismc_hmain0_s0_hrdata; 
wire            ismc_hmain0_s0_hready; 
wire    [1 :0]  ismc_hmain0_s0_hresp; 
wire            pmu_smc_hclk;         
wire            pmu_smc_hrst_b;       
wire    [31:0]  smc_hmain0_s2_hrdata; 
wire            smc_hmain0_s2_hready; 
wire    [1 :0]  smc_hmain0_s2_hresp;  
wire    [31:0]  smc_hmain0_s3_hrdata; 
wire            smc_hmain0_s3_hready; 
wire    [1 :0]  smc_hmain0_s3_hresp;  
wire    [31:0]  smc_hmain0_s4_hrdata; 
wire            smc_hmain0_s4_hready; 
wire    [1 :0]  smc_hmain0_s4_hresp;  

wire    [31:0]  hmain0_dummy3_s11_haddr;    
wire    [3 :0]  hmain0_dummy3_s11_hprot;    
wire            hmain0_dummy3_s11_hsel;     
wire    [2 :0]  hmain0_dummy3_s11_hsize;    
wire    [1 :0]  hmain0_dummy3_s11_htrans;   
wire    [31:0]  hmain0_dummy3_s11_hwdata;   
wire            hmain0_dummy3_s11_hwrite; 
wire    [31:0]  hmain0_dummy0_s7_haddr;     
wire    [3 :0]  hmain0_dummy0_s7_hprot;     
wire            hmain0_dummy0_s7_hsel;      
wire    [2 :0]  hmain0_dummy0_s7_hsize;     
wire    [1 :0]  hmain0_dummy0_s7_htrans;    
wire    [31:0]  hmain0_dummy0_s7_hwdata;    
wire            hmain0_dummy0_s7_hwrite;    
wire    [31:0]  hmain0_dummy1_s8_haddr;       
wire    [3 :0]  hmain0_dummy1_s8_hprot;     
wire            hmain0_dummy1_s8_hsel;      
wire    [2 :0]  hmain0_dummy1_s8_hsize;     
wire    [1 :0]  hmain0_dummy1_s8_htrans;    
wire    [31:0]  hmain0_dummy1_s8_hwdata;    
wire            hmain0_dummy1_s8_hwrite;    
wire    [31:0]  hmain0_dummy2_s9_haddr;       
wire    [3 :0]  hmain0_dummy2_s9_hprot;     
wire            hmain0_dummy2_s9_hsel;      
wire    [2 :0]  hmain0_dummy2_s9_hsize;     
wire    [1 :0]  hmain0_dummy2_s9_htrans;    
wire    [31:0]  hmain0_dummy2_s9_hwdata;    
wire            hmain0_dummy2_s9_hwrite; 

wire    [31:0]  dummy0_hmain0_s7_hrdata;    
wire            dummy0_hmain0_s7_hready;    
wire    [1 :0]  dummy0_hmain0_s7_hresp;     
wire    [31:0]  dummy1_hmain0_s8_hrdata;    
wire            dummy1_hmain0_s8_hready;    
wire    [1 :0]  dummy1_hmain0_s8_hresp;     
wire    [31:0]  dummy2_hmain0_s9_hrdata;    
wire            dummy2_hmain0_s9_hready;    
wire    [1 :0]  dummy2_hmain0_s9_hresp;     
wire    [31:0]  dummy3_hmain0_s11_hrdata;   
wire            dummy3_hmain0_s11_hready;   
wire    [1 :0]  dummy3_hmain0_s11_hresp; 

smu_top  x_smu1_top (
  .hmain0_ismc_s0_haddr  (hmain0_ismc_s0_haddr ),
  .hmain0_ismc_s0_hprot  (hmain0_ismc_s0_hprot ),
  .hmain0_ismc_s0_hsel   (hmain0_ismc_s0_hsel  ),
  .hmain0_ismc_s0_hsize  (hmain0_ismc_s0_hsize ),
  .hmain0_ismc_s0_htrans (hmain0_ismc_s0_htrans),
  .hmain0_ismc_s0_hwdata (hmain0_ismc_s0_hwdata),
  .hmain0_ismc_s0_hwrite (hmain0_ismc_s0_hwrite),
  .hmain0_smc_s2_haddr   (hmain0_smc_s2_haddr  ),
  .hmain0_smc_s2_hprot   (hmain0_smc_s2_hprot  ),
  .hmain0_smc_s2_hsel    (hmain0_smc_s2_hsel   ),
  .hmain0_smc_s2_hsize   (hmain0_smc_s2_hsize  ),
  .hmain0_smc_s2_htrans  (hmain0_smc_s2_htrans ),
  .hmain0_smc_s2_hwdata  (hmain0_smc_s2_hwdata ),
  .hmain0_smc_s2_hwrite  (hmain0_smc_s2_hwrite ),
  .hmain0_smc_s3_haddr   (hmain0_smc_s3_haddr  ),
  .hmain0_smc_s3_hprot   (hmain0_smc_s3_hprot  ),
  .hmain0_smc_s3_hsel    (hmain0_smc_s3_hsel   ),
  .hmain0_smc_s3_hsize   (hmain0_smc_s3_hsize  ),
  .hmain0_smc_s3_htrans  (hmain0_smc_s3_htrans ),
  .hmain0_smc_s3_hwdata  (hmain0_smc_s3_hwdata ),
  .hmain0_smc_s3_hwrite  (hmain0_smc_s3_hwrite ),
  .hmain0_smc_s4_haddr   (hmain0_smc_s4_haddr  ),
  .hmain0_smc_s4_hprot   (hmain0_smc_s4_hprot  ),
  .hmain0_smc_s4_hsel    (hmain0_smc_s4_hsel   ),
  .hmain0_smc_s4_hsize   (hmain0_smc_s4_hsize  ),
  .hmain0_smc_s4_htrans  (hmain0_smc_s4_htrans ),
  .hmain0_smc_s4_hwdata  (hmain0_smc_s4_hwdata ),
  .hmain0_smc_s4_hwrite  (hmain0_smc_s4_hwrite ),

  //TODO:1111
  .hmain0_imemdummy0_s1_haddr   (hmain0_imemdummy0_s1_haddr  ),
  .hmain0_imemdummy0_s1_hprot   (hmain0_imemdummy0_s1_hprot  ),
  .hmain0_imemdummy0_s1_hsel    (hmain0_imemdummy0_s1_hsel   ),
  .hmain0_imemdummy0_s1_hsize   (hmain0_imemdummy0_s1_hsize  ),
  .hmain0_imemdummy0_s1_htrans  (hmain0_imemdummy0_s1_htrans ),
  .hmain0_imemdummy0_s1_hwdata  (hmain0_imemdummy0_s1_hwdata ),
  .hmain0_imemdummy0_s1_hwrite  (hmain0_imemdummy0_s1_hwrite ),

  .hmain0_dummy3_s11_haddr (hmain0_dummy3_s11_haddr ),    
  .hmain0_dummy3_s11_hprot (hmain0_dummy3_s11_hprot ),    
  .hmain0_dummy3_s11_hsel  (hmain0_dummy3_s11_hsel  ),     
  .hmain0_dummy3_s11_hsize (hmain0_dummy3_s11_hsize ),    
  .hmain0_dummy3_s11_htrans(hmain0_dummy3_s11_htrans),   
  .hmain0_dummy3_s11_hwdata(hmain0_dummy3_s11_hwdata),   
  .hmain0_dummy3_s11_hwrite(hmain0_dummy3_s11_hwrite), 
  .hmain0_dummy0_s7_haddr  (hmain0_dummy0_s7_haddr  ),     
  .hmain0_dummy0_s7_hprot  (hmain0_dummy0_s7_hprot  ),     
  .hmain0_dummy0_s7_hsel   (hmain0_dummy0_s7_hsel   ),      
  .hmain0_dummy0_s7_hsize  (hmain0_dummy0_s7_hsize  ),     
  .hmain0_dummy0_s7_htrans (hmain0_dummy0_s7_htrans ),    
  .hmain0_dummy0_s7_hwdata (hmain0_dummy0_s7_hwdata ),    
  .hmain0_dummy0_s7_hwrite (hmain0_dummy0_s7_hwrite ),    
  .hmain0_dummy1_s8_haddr  (/*hmain0_dummy1_s8_haddr  */),       
  .hmain0_dummy1_s8_hprot  (/*hmain0_dummy1_s8_hprot  */),     
  .hmain0_dummy1_s8_hsel   (/*hmain0_dummy1_s8_hsel   */),      
  .hmain0_dummy1_s8_hsize  (/*hmain0_dummy1_s8_hsize  */),     
  .hmain0_dummy1_s8_htrans (/*hmain0_dummy1_s8_htrans */),    
  .hmain0_dummy1_s8_hwdata (/*hmain0_dummy1_s8_hwdata */),    
  .hmain0_dummy1_s8_hwrite (/*hmain0_dummy1_s8_hwrite */),    
  .hmain0_dummy2_s9_haddr  (/*hmain0_dummy2_s9_haddr  */),       
  .hmain0_dummy2_s9_hprot  (/*hmain0_dummy2_s9_hprot  */),     
  .hmain0_dummy2_s9_hsel   (/*hmain0_dummy2_s9_hsel   */),      
  .hmain0_dummy2_s9_hsize  (/*hmain0_dummy2_s9_hsize  */),     
  .hmain0_dummy2_s9_htrans (/*hmain0_dummy2_s9_htrans */),    
  .hmain0_dummy2_s9_hwdata (/*hmain0_dummy2_s9_hwdata */),    
  .hmain0_dummy2_s9_hwrite (/*hmain0_dummy2_s9_hwrite */), 

  .ismc_hmain0_s0_hrdata (ismc_hmain0_s0_hrdata),
  .ismc_hmain0_s0_hready (ismc_hmain0_s0_hready),
  .ismc_hmain0_s0_hresp  (ismc_hmain0_s0_hresp ),
  .pmu_smc_hclk          (pmu_smc_hclk         ),
  .pmu_smc_hrst_b        (pmu_smc_hrst_b       ),
  .smc_hmain0_s2_hrdata  (smc_hmain0_s2_hrdata ),
  .smc_hmain0_s2_hready  (smc_hmain0_s2_hready ),
  .smc_hmain0_s2_hresp   (smc_hmain0_s2_hresp  ),
  .smc_hmain0_s3_hrdata  (smc_hmain0_s3_hrdata ),
  .smc_hmain0_s3_hready  (smc_hmain0_s3_hready ),
  .smc_hmain0_s3_hresp   (smc_hmain0_s3_hresp  ),
  .smc_hmain0_s4_hrdata  (smc_hmain0_s4_hrdata ),
  .smc_hmain0_s4_hready  (smc_hmain0_s4_hready ),
  .smc_hmain0_s4_hresp   (smc_hmain0_s4_hresp  ),

  .imemdummy0_hmain0_s1_hrdata  (imemdummy0_hmain0_s1_hrdata),
  .imemdummy0_hmain0_s1_hready  (imemdummy0_hmain0_s1_hready),
  .imemdummy0_hmain0_s1_hresp   (imemdummy0_hmain0_s1_hresp),

  .dummy0_hmain0_s7_hrdata  (dummy0_hmain0_s7_hrdata ),    
  .dummy0_hmain0_s7_hready  (dummy0_hmain0_s7_hready ),    
  .dummy0_hmain0_s7_hresp   (dummy0_hmain0_s7_hresp  ),     
  .dummy1_hmain0_s8_hrdata  (dummy1_hmain0_s8_hrdata ),    
  .dummy1_hmain0_s8_hready  (dummy1_hmain0_s8_hready ),    
  .dummy1_hmain0_s8_hresp   (dummy1_hmain0_s8_hresp  ),     
  .dummy2_hmain0_s9_hrdata  (dummy2_hmain0_s9_hrdata ),    
  .dummy2_hmain0_s9_hready  (dummy2_hmain0_s9_hready ),    
  .dummy2_hmain0_s9_hresp   (dummy2_hmain0_s9_hresp  ),     
  .dummy3_hmain0_s11_hrdata (dummy3_hmain0_s11_hrdata),   
  .dummy3_hmain0_s11_hready (dummy3_hmain0_s11_hready),   
  .dummy3_hmain0_s11_hresp  (dummy3_hmain0_s11_hresp )

);


endmodule
